module sbox_aes (
    input  [7:0] X,   // 8-bit input
    output reg [7:0] Y  // 8-bit output
);

always @(*) begin
    case (X)
        8'b00000000: Y = 8'b01100011;  // '63'
        8'b00000001: Y = 8'b01111100;  // '7c'
        8'b00000010: Y = 8'b01110111;  // '77'
        8'b00000011: Y = 8'b01111011;  // '7b'
        8'b00000100: Y = 8'b11110010;  // 'f2'
        8'b00000101: Y = 8'b01101011;  // '6b'
        8'b00000110: Y = 8'b01101111;  // '6f'
        8'b00000111: Y = 8'b11000101;  // 'c5'
        8'b00001000: Y = 8'b00110000;  // '30'
        8'b00001001: Y = 8'b00000001;  // '01'
        8'b00001010: Y = 8'b01100111;  // '67'
        8'b00001011: Y = 8'b00101011;  // '2b'
        8'b00001100: Y = 8'b11111110;  // 'fe'
        8'b00001101: Y = 8'b11010111;  // 'd7'
        8'b00001110: Y = 8'b10101011;  // 'ab'
        8'b00001111: Y = 8'b01110110;  // '76'
        8'b00010000: Y = 8'b11001010;  // 'ca'
        8'b00010001: Y = 8'b10000010;  // '82'
        8'b00010010: Y = 8'b11001001;  // 'c9'
        8'b00010011: Y = 8'b01111101;  // '7d'
        8'b00010100: Y = 8'b11111010;  // 'fa'
        8'b00010101: Y = 8'b01011001;  // '59'
        8'b00010110: Y = 8'b01000111;  // '47'
        8'b00010111: Y = 8'b11110000;  // 'f0'
        8'b00011000: Y = 8'b10101101;  // 'ad'
        8'b00011001: Y = 8'b11010100;  // 'd4'
        8'b00011010: Y = 8'b10100010;  // 'a2'
        8'b00011011: Y = 8'b10101111;  // 'af'
        8'b00011100: Y = 8'b10011100;  // '9c'
        8'b00011101: Y = 8'b10100100;  // 'a4'
        8'b00011110: Y = 8'b01110010;  // '72'
        8'b00011111: Y = 8'b11000000;  // 'c0'
        8'b00100000: Y = 8'b10110111;  // 'b7'
        8'b00100001: Y = 8'b11111101;  // 'fd'
        8'b00100010: Y = 8'b10010011;  // '93'
        8'b00100011: Y = 8'b00100110;  // '26'
        8'b00100100: Y = 8'b00110110;  // '36'
        8'b00100101: Y = 8'b00111111;  // '3f'
        8'b00100110: Y = 8'b11110111;  // 'f7'
        8'b00100111: Y = 8'b11001100;  // 'cc'
        8'b00101000: Y = 8'b00110100;  // '34'
        8'b00101001: Y = 8'b10100101;  // 'a5'
        8'b00101010: Y = 8'b11100101;  // 'e5'
        8'b00101011: Y = 8'b11110001;  // 'f1'
        8'b00101100: Y = 8'b01110001;  // '71'
        8'b00101101: Y = 8'b11011000;  // 'd8'
        8'b00101110: Y = 8'b00110001;  // '31'
        8'b00101111: Y = 8'b00010101;  // '15'
        8'b00110000: Y = 8'b00000100;  // '04'
        8'b00110001: Y = 8'b11000111;  // 'c7'
        8'b00110010: Y = 8'b00100011;  // '23'
        8'b00110011: Y = 8'b11000011;  // 'c3'
        8'b00110100: Y = 8'b00011000;  // '18'
        8'b00110101: Y = 8'b10010110;  // '96'
        8'b00110110: Y = 8'b00000101;  // '05'
        8'b00110111: Y = 8'b10011010;  // '9a'
        8'b00111000: Y = 8'b00000111;  // '07'
        8'b00111001: Y = 8'b00010010;  // '12'
        8'b00111010: Y = 8'b10000000;  // '80'
        8'b00111011: Y = 8'b11100010;  // 'e2'
        8'b00111100: Y = 8'b11101011;  // 'eb'
        8'b00111101: Y = 8'b00100111;  // '27'
        8'b00111110: Y = 8'b10110010;  // 'b2'
        8'b00111111: Y = 8'b01110101;  // '75'
        8'b01000000: Y = 8'b00001001;  // '09'
        8'b01000001: Y = 8'b10000011;  // '83'
        8'b01000010: Y = 8'b00101100;  // '2c'
        8'b01000011: Y = 8'b00011010;  // '1a'
        8'b01000100: Y = 8'b00011011;  // '1b'
        8'b01000101: Y = 8'b01101110;  // '6e'
        8'b01000110: Y = 8'b01011010;  // '5a'
        8'b01000111: Y = 8'b10100000;  // 'a0'
        8'b01001000: Y = 8'b01010010;  // '52'
        8'b01001001: Y = 8'b00111011;  // '3b'
        8'b01001010: Y = 8'b11010110;  // 'd6'
        8'b01001011: Y = 8'b10110011;  // 'b3'
        8'b01001100: Y = 8'b00101001;  // '29'
        8'b01001101: Y = 8'b11100011;  // 'e3'
        8'b01001110: Y = 8'b00101111;  // '2f'
        8'b01001111: Y = 8'b10000100;  // '84'
        8'b01010000: Y = 8'b01010011;  // '53'
        8'b01010001: Y = 8'b11010001;  // 'd1'
        8'b01010010: Y = 8'b00000000;  // '00'
        8'b01010011: Y = 8'b11101101;  // 'ed'
        8'b01010100: Y = 8'b00100000;  // '20'
        8'b01010101: Y = 8'b11111100;  // 'fc'
        8'b01010110: Y = 8'b10110001;  // 'b1'
        8'b01010111: Y = 8'b01011011;  // '5b'
        8'b01011000: Y = 8'b01101010;  // '6a'
        8'b01011001: Y = 8'b11001011;  // 'cb'
        8'b01011010: Y = 8'b10111110;  // 'be'
        8'b01011011: Y = 8'b00111001;  // '39'
        8'b01011100: Y = 8'b01001010;  // '4a'
        8'b01011101: Y = 8'b01001100;  // '4c'
        8'b01011110: Y = 8'b01011000;  // '58'
        8'b01011111: Y = 8'b11001111;  // 'cf'
        8'b01100000: Y = 8'b11010000;  // 'd0'
        8'b01100001: Y = 8'b11101111;  // 'ef'
        8'b01100010: Y = 8'b10101010;  // 'aa'
        8'b01100011: Y = 8'b11111011;  // 'fb'
        8'b01100100: Y = 8'b01000011;  // '43'
        8'b01100101: Y = 8'b01001101;  // '4d'
        8'b01100110: Y = 8'b00110011;  // '33'
        8'b01100111: Y = 8'b10000101;  // '85'
        8'b01101000: Y = 8'b01000101;  // '45'
        8'b01101001: Y = 8'b11111001;  // 'f9'
        8'b01101010: Y = 8'b00000010;  // '02'
        8'b01101011: Y = 8'b01111111;  // '7f'
        8'b01101100: Y = 8'b01010000;  // '50'
        8'b01101101: Y = 8'b00111100;  // '3c'
        8'b01101110: Y = 8'b10011111;  // '9f'
        8'b01101111: Y = 8'b10101000;  // 'a8'
        8'b01110000: Y = 8'b01010001;  // '51'
        8'b01110001: Y = 8'b10100011;  // 'a3'
        8'b01110010: Y = 8'b01000000;  // '40'
        8'b01110011: Y = 8'b10001111;  // '8f'
        8'b01110100: Y = 8'b10010010;  // '92'
        8'b01110101: Y = 8'b10011101;  // '9d'
        8'b01110110: Y = 8'b00111000;  // '38'
        8'b01110111: Y = 8'b11110101;  // 'f5'
        8'b01111000: Y = 8'b10111100;  // 'bc'
        8'b01111001: Y = 8'b10110110;  // 'b6'
        8'b01111010: Y = 8'b11011010;  // 'da'
        8'b01111011: Y = 8'b00100001;  // '21'
        8'b01111100: Y = 8'b00010000;  // '10'
        8'b01111101: Y = 8'b11111111;  // 'ff'
        8'b01111110: Y = 8'b11110011;  // 'f3'
        8'b01111111: Y = 8'b11010010;  // 'd2'
        8'b10000000: Y = 8'b11001101;  // 'cd'
        8'b10000001: Y = 8'b00001100;  // '0c'
        8'b10000010: Y = 8'b00010011;  // '13'
        8'b10000011: Y = 8'b11101100;  // 'ec'
        8'b10000100: Y = 8'b01011111;  // '5f'
        8'b10000101: Y = 8'b10010111;  // '97'
        8'b10000110: Y = 8'b01000100;  // '44'
        8'b10000111: Y = 8'b00010111;  // '17'
        8'b10001000: Y = 8'b11000100;  // 'c4'
        8'b10001001: Y = 8'b10100111;  // 'a7'
        8'b10001010: Y = 8'b01111110;  // '7e'
        8'b10001011: Y = 8'b00111101;  // '3d'
        8'b10001100: Y = 8'b01100100;  // '64'
        8'b10001101: Y = 8'b01011101;  // '5d'
        8'b10001110: Y = 8'b00011001;  // '19'
        8'b10001111: Y = 8'b01110011;  // '73'
        8'b10010000: Y = 8'b01100000;  // '60'
        8'b10010001: Y = 8'b10000001;  // '81'
        8'b10010010: Y = 8'b01001111;  // '4f'
        8'b10010011: Y = 8'b11011100;  // 'dc'
        8'b10010100: Y = 8'b00100010;  // '22'
        8'b10010101: Y = 8'b00101010;  // '2a'
        8'b10010110: Y = 8'b10010000;  // '90'
        8'b10010111: Y = 8'b10001000;  // '88'
        8'b10011000: Y = 8'b01000110;  // '46'
        8'b10011001: Y = 8'b11101110;  // 'ee'
        8'b10011010: Y = 8'b10111000;  // 'b8'
        8'b10011011: Y = 8'b00010100;  // '14'
        8'b10011100: Y = 8'b11011110;  // 'de'
        8'b10011101: Y = 8'b01011110;  // '5e'
        8'b10011110: Y = 8'b00001011;  // '0b'
        8'b10011111: Y = 8'b11011011;  // 'db'
        8'b10100000: Y = 8'b11100000;  // 'e0'
        8'b10100001: Y = 8'b00110010;  // '32'
        8'b10100010: Y = 8'b00111010;  // '3a'
        8'b10100011: Y = 8'b00001010;  // '0a'
        8'b10100100: Y = 8'b01001001;  // '49'
        8'b10100101: Y = 8'b00000110;  // '06'
        8'b10100110: Y = 8'b00100100;  // '24'
        8'b10100111: Y = 8'b01011100;  // '5c'
        8'b10101000: Y = 8'b11000010;  // 'c2'
        8'b10101001: Y = 8'b11010011;  // 'd3'
        8'b10101010: Y = 8'b10101100;  // 'ac'
        8'b10101011: Y = 8'b01100010;  // '62'
        8'b10101100: Y = 8'b10010001;  // '91'
        8'b10101101: Y = 8'b10010101;  // '95'
        8'b10101110: Y = 8'b11100100;  // 'e4'
        8'b10101111: Y = 8'b01111001;  // '79'
        8'b10110000: Y = 8'b11100111;  // 'e7'
        8'b10110001: Y = 8'b11001000;  // 'c8'
        8'b10110010: Y = 8'b00110111;  // '37'
        8'b10110011: Y = 8'b01101101;  // '6d'
        8'b10110100: Y = 8'b10001101;  // '8d'
        8'b10110101: Y = 8'b11010101;  // 'd5'
        8'b10110110: Y = 8'b01001110;  // '4e'
        8'b10110111: Y = 8'b10101001;  // 'a9'
        8'b10111000: Y = 8'b01101100;  // '6c'
        8'b10111001: Y = 8'b01010110;  // '56'
        8'b10111010: Y = 8'b11110100;  // 'f4'
        8'b10111011: Y = 8'b11101010;  // 'ea'
        8'b10111100: Y = 8'b01100101;  // '65'
        8'b10111101: Y = 8'b01111010;  // '7a'
        8'b10111110: Y = 8'b10101110;  // 'ae'
        8'b10111111: Y = 8'b00001000;  // '08'
        8'b11000000: Y = 8'b10111010;  // 'ba'
        8'b11000001: Y = 8'b01111000;  // '78'
        8'b11000010: Y = 8'b00100101;  // '25'
        8'b11000011: Y = 8'b00101110;  // '2e'
        8'b11000100: Y = 8'b00011100;  // '1c'
        8'b11000101: Y = 8'b10100110;  // 'a6'
        8'b11000110: Y = 8'b10110100;  // 'b4'
        8'b11000111: Y = 8'b11000110;  // 'c6'
        8'b11001000: Y = 8'b11101000;  // 'e8'
        8'b11001001: Y = 8'b11011101;  // 'dd'
        8'b11001010: Y = 8'b01110100;  // '74'
        8'b11001011: Y = 8'b00011111;  // '1f'
        8'b11001100: Y = 8'b01001011;  // '4b'
        8'b11001101: Y = 8'b10111101;  // 'bd'
        8'b11001110: Y = 8'b10001011;  // '8b'
        8'b11001111: Y = 8'b10001010;  // '8a'
        8'b11010000: Y = 8'b01110000;  // '70'
        8'b11010001: Y = 8'b00111110;  // '3e'
        8'b11010010: Y = 8'b10110101;  // 'b5'
        8'b11010011: Y = 8'b01100110;  // '66'
        8'b11010100: Y = 8'b01001000;  // '48'
        8'b11010101: Y = 8'b00000011;  // '03'
        8'b11010110: Y = 8'b11110110;  // 'f6'
        8'b11010111: Y = 8'b00001110;  // '0e'
        8'b11011000: Y = 8'b01100001;  // '61'
        8'b11011001: Y = 8'b00110101;  // '35'
        8'b11011010: Y = 8'b01010111;  // '57'
        8'b11011011: Y = 8'b10111001;  // 'b9'
        8'b11011100: Y = 8'b10000110;  // '86'
        8'b11011101: Y = 8'b11000001;  // 'c1'
        8'b11011110: Y = 8'b00011101;  // '1d'
        8'b11011111: Y = 8'b10011110;  // '9e'
        8'b11100000: Y = 8'b11100001;  // 'e1'
        8'b11100001: Y = 8'b11111000;  // 'f8'
        8'b11100010: Y = 8'b10011000;  // '98'
        8'b11100011: Y = 8'b00010001;  // '11'
        8'b11100100: Y = 8'b01101001;  // '69'
        8'b11100101: Y = 8'b11011001;  // 'd9'
        8'b11100110: Y = 8'b10001110;  // '8e'
        8'b11100111: Y = 8'b10010100;  // '94'
        8'b11101000: Y = 8'b10011011;  // '9b'
        8'b11101001: Y = 8'b00011110;  // '1e'
        8'b11101010: Y = 8'b10000111;  // '87'
        8'b11101011: Y = 8'b11101001;  // 'e9'
        8'b11101100: Y = 8'b11001110;  // 'ce'
        8'b11101101: Y = 8'b01010101;  // '55'
        8'b11101110: Y = 8'b00101000;  // '28'
        8'b11101111: Y = 8'b11011111;  // 'df'
        8'b11110000: Y = 8'b10001100;  // '8c'
        8'b11110001: Y = 8'b10100001;  // 'a1'
        8'b11110010: Y = 8'b10001001;  // '89'
        8'b11110011: Y = 8'b00001101;  // '0d'
        8'b11110100: Y = 8'b10111111;  // 'bf'
        8'b11110101: Y = 8'b11100110;  // 'e6'
        8'b11110110: Y = 8'b01000010;  // '42'
        8'b11110111: Y = 8'b01101000;  // '68'
        8'b11111000: Y = 8'b01000001;  // '41'
        8'b11111001: Y = 8'b10011001;  // '99'
        8'b11111010: Y = 8'b00101101;  // '2d'
        8'b11111011: Y = 8'b00001111;  // '0f'
        8'b11111100: Y = 8'b10110000;  // 'b0'
        8'b11111101: Y = 8'b01010100;  // '54'
        8'b11111110: Y = 8'b10111011;  // 'bb'
        8'b11111111: Y = 8'b00010110;  // '16'
    endcase
end


endmodule
